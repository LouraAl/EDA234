----------------------------------------------------------------------------------                         
-- Company:                                                                                                
-- Engineer:                                                                                               
--                                                                                                         
-- Create Date: 11/06/2025 02:25:02 PM                                                                     
-- Design Name:                                                                                            
-- Module Name: demo - Behavioral                                                                          
-- Project Name:                                                                                           
-- Target Devices:                                                                                         
-- Tool Versions:                                                                                          
-- Description:                                                                                            
--                                                                                                         
-- Dependencies:                                                                                           
--                                                                                                         
-- Revision:                                                                                               
-- Revision 0.01 - File Created                                                                            
-- Additional Comments:                                                                                    
--                                                                                                         
----------------------------------------------------------------------------------                         
                                                                                                           
                                                                                                           
library IEEE;                                                                                              
use IEEE.STD_LOGIC_1164.ALL;                                                                               
                                                                                                           
-- Uncomment the following library declaration if using                                                    
-- arithmetic functions with Signed or Unsigned values                                                     
use IEEE.NUMERIC_STD.ALL;
                                                                                
                                                                                                           
-- Uncomment the following library declaration if instantiating                                            
-- any Xilinx leaf cells in this code.                                                                     
--library UNISIM;                                                                                          
--use UNISIM.VComponents.all;                                                                              
                                                                                                           
entity LAB1H1 is     
  generic( 
	constant  CTRL_max :  natural := 25 - 1; --refresh per 200Hz (250 000) on the displays or 25 for simulation                                        
  	constant sec_pulse_max :natural := 1000 - 1); --refresh per 1Hz (100 000 000) for 1 second counter, or 1000 for simulation
	                                                                                       
  port ( CLK: in std_logic;
	 RESET: in std_logic;                                                                                                                                      
         SEG: out std_logic_vector(7 downto 0);                                                          
         AN : out STD_LOGIC_VECTOR (7 downto 0));                                                        
end LAB1H1;                                                                                                 
                                                                                                           
architecture Behavioral of LAB1H1 is 
  signal one_digit   : unsigned(3 downto 0);  -- selects digit 0..9
  signal ten_digit    : unsigned(3 downto 0);  -- selects digit 0..9 
  
  signal sec_cnt   : unsigned(3 downto 0);  -- enough for 9 second count
  signal ten_sec_cnt   : unsigned(3 downto 0);  -- enough for 50 second count
  signal mux_select : std_logic; 

  signal seg_pat10  : std_logic_vector(7 downto 0);
  signal seg_pat1 : std_logic_vector(7 downto 0);                                                                                                                                                                                                                                                                                                                                                                                                              
 
 Begin 
COUNTER: PROCESS(CLK, reset) 

   variable CTRL : unsigned(18 downto 0);
   variable sec_pulse : unsigned(27 downto 0);
  Begin
    if reset = '1' then
	  ten_sec_cnt <= (others => '0');
	  sec_pulse := (others => '0');
	  sec_cnt <= (others => '0');
	  mux_select <= '0';
	  CTRL := (others => '0');

    elsif rising_edge(CLK) then
	  if sec_pulse = sec_pulse_max then
		sec_pulse := (others => '0');
		if sec_cnt = 9 then 
		   sec_cnt <= (others => '0');
		   ten_sec_cnt <= ten_sec_cnt + 1;
			if ten_sec_cnt = 5 then 
		   	ten_sec_cnt <= (others => '0');
			end if;
		else
		   sec_cnt <= sec_cnt + 1;
		end if; 
	  else 
		sec_pulse := sec_pulse + 1;
	  end if;
	  
	  if CTRL = CTRL_max then
		CTRL := (others => '0');
		mux_select <= not mux_select;
	  else
		CTRL := CTRL + 1;
	  end if;
    end if;
END PROCESS COUNTER;


SecToBits: PROCESS (sec_cnt)  
  Begin
      ten_digit <= ten_sec_cnt;
      one_digit <= sec_cnt;
END PROCESS SecToBits;
  
DISPLAY: PROCESS (ten_digit, one_digit)
  Begin                                                                                                  
   	CASE one_digit IS
				WHEN "0000" =>
					seg_pat1 <="11000000"; --0
				WHEN "0001" =>
					seg_pat1 <="11111001"; --1
				WHEN "0010" =>
					seg_pat1 <="10100100"; --2
				WHEN "0011" =>
					seg_pat1 <="10110000"; --3
				WHEN "0100" =>
					seg_pat1 <="10011001"; --4
				WHEN "0101" =>
					seg_pat1 <="10010010"; --5
				WHEN "0110" =>
					seg_pat1 <="10000010"; --6
				WHEN "0111" =>
					seg_pat1 <="11111000"; --7
				WHEN "1000" =>
					seg_pat1 <="10000000"; --8
				WHEN "1001" =>
					seg_pat1 <="10010000"; --9
				WHEN others =>
					seg_pat1 <="11111111"; --off
	END CASE;
	CASE ten_digit IS
				WHEN "0000" =>
					seg_pat10 <="11000000"; --0
				WHEN "0001" =>
					seg_pat10 <="11111001"; --1
				WHEN "0010" =>
					seg_pat10 <="10100100"; --2
				WHEN "0011" =>
					seg_pat10 <="10110000"; --3
				WHEN "0100" =>
					seg_pat10 <="10011001"; --4
				WHEN "0101" =>
					seg_pat10 <="10010010"; --5
				WHEN "0110" =>
					seg_pat10 <="10000010"; --6
				WHEN "0111" =>
					seg_pat10 <="11111000"; --7
				WHEN "1000" =>
					seg_pat10 <="10000000"; --8
				WHEN "1001" =>
					seg_pat10 <="10010000"; --9
				WHEN others =>
					seg_pat10 <="11111111"; --off
	END CASE; --SW
END PROCESS DISPLAY;   

OUTPUT_DISPLAY: PROCESS (mux_select, seg_pat10, seg_pat1)
    Begin 
	if mux_select = '0' then 
	   AN (7 downto 0) <= "11111110";
	   Seg <= seg_pat1(7 downto 0);
	else 
	   AN (7 downto 0) <= "11111101"; 
	   Seg <= seg_pat10(7 downto 0);
	end if; 
END PROCESS OUTPUT_DISPLAY;                                                                                                     
                                                                            
end Behavioral;                                                
